
module if_if_stages_tb (
    
);
    
endmodule